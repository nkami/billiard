


module	back_ground	(	

					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0]	pixelX,
					input logic	[10:0]	pixelY,
					input logic menu_state, // game menu is currently open
					input logic game_state, // game is currently running
					input logic end_state,  // game ended
					input logic win,  // game won

					output logic [7:0]	BG_RGB
);

// maybe for testing we should use them with LPM_CONST
parameter int	topLeftTableX = 60;
parameter int	topLeftTableY = 90;
parameter int	tableWidth = 520;
parameter int	tableHeight = 270;
parameter int	woodWidth = 20;
parameter int  topLeftMenuX = 150;
parameter int  topLeftMenuY = 150;
parameter int  topLeftWinX = 150;
parameter int  topLeftWinY = 175;
parameter int  topLeftLoseX = 150;
parameter int  topLeftLoseY = 175;
parameter int  topLeftStrikesX = 285;
parameter int  topLeftStrikesY = 0;


// the holes are numbered from 1 to 6 clockwise starting from the upper left hole
const int	topLeftHole1X = 65;
const int	topLeftHole1Y = 95;

const int	topLeftHole2X = 300;
const int	topLeftHole2Y = 95;

const int	topLeftHole3X = 543;
const int	topLeftHole3Y = 95;

const int	topLeftHole4X = 543;
const int	topLeftHole4Y = 322;

const int	topLeftHole5X = 300;
const int	topLeftHole5Y = 322;

const int	topLeftHole6X = 65;
const int	topLeftHole6Y = 322;

// bitmaps for table holes, menu text, winning text and losing text

localparam  int HOLE_WIDTH_X = 32;
localparam  int HOLE_HEIGHT_Y = 32;

logic [0:HOLE_HEIGHT_Y-1] [0:HOLE_WIDTH_X-1] [1-1:0] hole_colors = {
{1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, },
{1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, },
{1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, },
{1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, },
{1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, },
{1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, },
{1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, },
{1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, },
{1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, },
{1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, },
{1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, },
{1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, },
{1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, },
{1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, },
{1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, },
{1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, },
{1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, },
{1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, },
{1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, },
{1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, },
{1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, },
{1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, },
{1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, },
{1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, },
{1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, },
{1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, },
{1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, },
{1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, },
{1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, },
{1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, },
{1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, },
{1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, }
};


localparam  int MENU_WIDTH_X = 350;
localparam  int MENU_HEIGHT_Y = 100;

logic [0:MENU_HEIGHT_Y-1] [1*MENU_WIDTH_X-1:0] menu_colors = {
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000011111000000000111111000000000001111110000001111111100000011111111111111111001111111111111111110000000000011111100011111111110000001111100011111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000001111000000000011111000000000001111100000000011111000000000111111111111110001111111111111111110000000000011111100011111111100000000011110001111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111000111001111110001111001111111111111000111110001110001111100011111111111100001111111111111111110011111111111111000001111111000111110001111001111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111100111001111111001111001111111111111001111111001110011111110011111111110000001111111111111111110011111111111111001001111111001111111001111000111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111100111001111111001111001111111111111001111111111110011111111111111111110011001111100111111111110011111111111111001001111111001111111111111100011000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111100111001111110001111001111111111111000111111111110001111111111111111111111001111100111111111110011111111111110011100111111000111111111111110011001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111000111000000000011111000000000011111100000011111111000000111111111111111111001111111111111111110000000000111110011100111111100000011111111110000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000001111000000000111111000000000011111111000000111111110000001111111111111111001111111111111111110000000000111100011100011111111000000111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000011111001110001111111001111111111111111111100011111111111000111111111111111001111111111111111110011111111111100000000011111111111100011111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111001111000111111001111111111111111111111001111111111110011111111111111001111111111111111110011111111111100000000011111111111111001111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111001111100111111001111111111110011111111001100111111110011111111111111001111111111111111110011111111111001111111001110011111111001111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111001111100011111001111111111110001111111001100011111110011111111111111001111111111111111110011111111111001111111001110001111111001111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111001111110001111001111111111111000111110001110001111100011111111111111001111111111111111110011111111111001111111001111000111110001111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111001111110001111000000000001111100000000011111000000000111111111111111001111100111111111110000000000010011111111100111100000000011111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111001111111000111000000000001111110000001111111100000011111111111111111001111100111111111110000000000010011111111100111110000001111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111110000000001111100000000011111100000000000111111000000111111110000001111111111111100000011111111111111110001111111110001110000000000011110000000001111110011100111111110011100011111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000111100000000001111100000000000111110000000001111100000000011111111111000000001111111111111110000111111100001110000000000011110000000000111110011100111111110011100001111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111110011111100011100111111000111100111111111111100011111000111000111110001111111110001111000111111111111110000111111100001110011111111111110011111100011110011100111111110011100001111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111110011111110011100111111100111100111111111111100111111100111001111111001111111110011111100111111111111110000111111100001110011111111111110011111110011110011100111111110011100001111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111110011111110011100111111100111100111111111111100111111111111001111111111111111111111111100110011111111110010011111001001110011111111111110011111110001110011100111111110011100100111110010011111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111110011111110011100111111000111100111111111111100011111111111000111111111111111111111111100110011111111110010011111001001110011111111111110011111111001110011100111111110011100100111110010011111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111110011111100011100000000001111100000000001111110000001111111100000011111111111111111111001111111111111110010011111001001110000000000111110011111111001110011100111111110011100100111110010011111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000111100000000011111100000000001111111100000011111111000000111111111111111110001111111111111110011001110011001110000000000111110011111111001110011100111111110011100110011100110011111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111110000000001111100111000111111100111111111111111111110001111111111100011111111111111110011111111111111110011001110011001110011111111111110011111111001110011100111111110011100110011100110011111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111100111100011111100111111111111111111111100111111111111001111111111111000111111111111111110011001110011001110011111111111110011111111001110011100111111110011100110011100110011111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111100111110011111100111111111111001111111100110011111111001111111111110001111111111111111110011100100111001110011111111111110011111110001110011100111111110011100111001001110011111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111100111110001111100111111111111000111111100110001111111001111111111100111111111111111111110011100100111001110011111111111110011111110011110011100011111100011100111001001110011111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111100111111000111100111111111111100011111000111000111110001111111111001111111111111111111110011100000111001110011111111111110011111100011110011110001111000111100111000001110011111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111100111111000111100000000000111110000000001111100000000011111111110000000000110011111111110011110001111001110000000000011110000000000111110011111000000001111100111100011110011111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111100111111100011100000000000111111000000111111110000001111111111110000000000110011111111110011110001111001110000000000011110000000011111110011111100000011111100111100011110011111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000001111100000000011111100000000000111111000000111111110000001111111111111100000111111111111111110011111111001111111000111111110000000001111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000111100000000001111100000000000111110000000001111100000000011111111111000000011111111111111110011111111001111111000111111110000000000111111000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111100011100111111000111100111111111111100011111000111000111110001111111110001110001111111111111110011111111001111110000011111110011111100011111001111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111110011100111111100111100111111111111100111111100111001111111001111111110011111001111111111111110011111111001111110010011111110011111110011111001111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111110011100111111100111100111111111111100111111111111001111111111111111111111111001110011111111110011111111001111110010011111110011111110011111001111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111110011100111111000111100111111111111100011111111111000111111111111111111111110011110011111111110011111111001111100111001111110011111100011111001111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111100011100000000001111100000000001111110000001111111100000011111111111111111000011111111111111110000000000001111100111001111110000000000111111001111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000111100000000011111100000000001111111100000011111111000000111111111111111000001111111111111110000000000001111000111000111110000000001111111001111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000001111100111000111111100111111111111111111110001111111111100011111111111111111000111111111111110011111111001111000000000111110011100011111111001111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111100111100011111100111111111111111111111100111111111111001111111111111111100111111111111110011111111001111000000000111110011110001111111001111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111100111110011111100111111111111001111111100110011111111001111111111111111100111111111111110011111111001110011111110011110011111001111111001111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111100111110001111100111111111111000111111100110001111111001111111110011111100111111111111110011111111001110011111110011110011111000111111001111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111100111111000111100111111111111100011111000111000111110001111111110001111001111111111111110011111111001110011111110011110011111100011111001111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111100111111000111100000000000111110000000001111100000000011111111111000000001110011111111110011111111001100111111111001110011111100011111000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111100111111100011100000000000111111000000111111110000001111111111111100000111110011111111110011111111001100111111111001110011111110001111000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{350'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111}
};



localparam  int WIN_WIDTH_X = 270;
localparam  int WIN_HEIGHT_Y = 70;

logic [0:WIN_HEIGHT_Y-1] [1*WIN_WIDTH_X-1:0] win_colors = {
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111100000111111111111111111000001111111111100000000011111111111111100001111111111111111100001111111111111111000011111111111110000000111111111111100001111111111100000000011111111111111000001111111111111111000011111111000011111111111111111111111111111},
{270'b111111111111111111111111110000011111111111111110000011111111110000000000000111111111111100001111111111111111100001111111111111111000001111111111110000000111111111111000001111111110000000000000111111111111000001111111111111111000011111111000011111111111111111111111111111},
{270'b111111111111111111111111111000011111111111111110000111111111000000000000000001111111111100001111111111111111100001111111111111111100001111111111110000000111111111111000011111111000000000000000001111111111000000111111111111111000011111111000011111111111111111111111111111},
{270'b111111111111111111111111111000001111111111111100000111111110000000000000000000111111111100001111111111111111100001111111111111111100001111111111100000000011111111111000011111110000000000000000000111111111000000011111111111111000011111111000011111111111111111111111111111},
{270'b111111111111111111111111111100000111111111111000001111111100000001111111000000011111111100001111111111111111100001111111111111111100001111111111100000000011111111111000011111100000001111111000000011111111000000011111111111111000011111111000011111111111111111111111111111},
{270'b111111111111111111111111111110000111111111111000011111111000000111111111110000001111111100001111111111111111100001111111111111111100001111111111100001000011111111111000011111000000111111111110000001111111000000001111111111111000011111111000011111111111111111111111111111},
{270'b111111111111111111111111111110000011111111110000011111110000001111111111111000000111111100001111111111111111100001111111111111111110000111111111100001000011111111110000111110000001111111111111000000111111000000000111111111111000011111111000011111111111111111111111111111},
{270'b111111111111111111111111111111000001111111100000111111110000011111111111111100000111111100001111111111111111100001111111111111111110000111111111000001000001111111110000111110000011111111111111100000111111000010000111111111111000011111111000011111111111111111111111111111},
{270'b111111111111111111111111111111100001111111100001111111100000111111111111111110000011111100001111111111111111100001111111111111111110000111111111000011100001111111110000111100000111111111111111110000011111000010000011111111111000011111111000011111111111111111111111111111},
{270'b111111111111111111111111111111100000111111000001111111100001111111111111111111000011111100001111111111111111100001111111111111111111000111111111000011100001111111110001111100001111111111111111111000011111000011000001111111111000011111111000011111111111111111111111111111},
{270'b111111111111111111111111111111110000011110000011111111100001111111111111111111000011111100001111111111111111100001111111111111111111000011111111000011100001111111100001111100001111111111111111111000011111000011100001111111111000011111111000011111111111111111111111111111},
{270'b111111111111111111111111111111111000011110000111111111000001111111111111111111000001111100001111111111111111100001111111111111111111000011111110000011100000111111100001111000001111111111111111111000001111000011100000111111111000011111111000011111111111111111111111111111},
{270'b111111111111111111111111111111111000001100000111111111000011111111111111111111100001111100001111111111111111100001111111111111111111000011111110000111110000111111100001111000011111111111111111111100001111000011110000011111111000011111111000011111111111111111111111111111},
{270'b111111111111111111111111111111111100000000001111111111000011111111111111111111100001111100001111111111111111100001111111111111111111100011111110000111110000111111100011111000011111111111111111111100001111000011111000011111111000011111111000011111111111111111111111111111},
{270'b111111111111111111111111111111111110000000011111111111000011111111111111111111100001111100001111111111111111100001111111111111111111100001111110000111110000111111000011111000011111111111111111111100001111000011111000001111111000011111111000011111111111111111111111111111},
{270'b111111111111111111111111111111111110000000011111111111000011111111111111111111100001111100001111111111111111100001111111111111111111100001111100001111111000011111000011111000011111111111111111111100001111000011111100000111111000011111111000011111111111111111111111111111},
{270'b111111111111111111111111111111111111000000111111111111000011111111111111111111100001111100001111111111111111100001111111111111111111100001111100001111111000011111000011111000011111111111111111111100001111000011111110000011111000011111111000011111111111111111111111111111},
{270'b111111111111111111111111111111111111100001111111111111000011111111111111111111100001111100001111111111111111100001111111111111111111110001111100001111111000011111000111111000011111111111111111111100001111000011111111000011111000011111111100111111111111111111111111111111},
{270'b111111111111111111111111111111111111100001111111111111000011111111111111111111100001111100001111111111111111100001111111111111111111110000111100001111111000011110000111111000011111111111111111111100001111000011111111000001111000011111111100111111111111111111111111111111},
{270'b111111111111111111111111111111111111100001111111111111000001111111111111111111000001111100001111111111111111100001111111111111111111110000111000011111111100001110000111111000001111111111111111111000001111000011111111100000111000011111111100111111111111111111111111111111},
{270'b111111111111111111111111111111111111100001111111111111100001111111111111111111000011111100001111111111111111100001111111111111111111111000111000011111111100001110001111111100001111111111111111111000011111000011111111110000111000011111111100111111111111111111111111111111},
{270'b111111111111111111111111111111111111100001111111111111100001111111111111111111000011111100001111111111111111100001111111111111111111111000111000011111111100001110001111111100001111111111111111111000011111000011111111110000011000011111111100111111111111111111111111111111},
{270'b111111111111111111111111111111111111100001111111111111100000111111111111111110000011111100000111111111111111000001111111111111111111111000011000011111111100001100001111111100000111111111111111110000011111000011111111111000001000011111111100111111111111111111111111111111},
{270'b111111111111111111111111111111111111100001111111111111110000011111111111111100000111111110000111111111111111000011111111111111111111111000010000111111111110000100001111111110000011111111111111100000111111000011111111111100001000011111111100111111111111111111111111111111},
{270'b111111111111111111111111111111111111100001111111111111110000001111111111111000000111111110000011111111111110000011111111111111111111111100010000111111111110000100011111111110000001111111111111000000111111000011111111111100000000011111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111100001111111111111111000000111111111110000001111111110000001111111111100000011111111111111111111111100010000111111111110000100011111111111000000111111111110000001111111000011111111111110000000011111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111100001111111111111111100000001111111000000011111111111000000011111110000000111111111111111111111111100000000111111111110000000011111111111100000001111111000000011111111000011111111111111000000011111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111100001111111111111111110000000000000000000111111111111100000000000000000001111111111111111111111111100000001111111111111000000011111111111110000000000000000000111111111000011111111111111000000011111111000011111111111111111111111111111},
{270'b111111111111111111111111111111111111100001111111111111111111000000000000000001111111111111110000000000000000011111111111111111111111111110000001111111111111000000111111111111111000000000000000001111111111000011111111111111100000011111111000011111111111111111111111111111},
{270'b111111111111111111111111111111111111100001111111111111111111110000000000000111111111111111111000000000000000111111111111111111111111111110000001111111111111000000111111111111111110000000000000111111111111000011111111111111110000011111111000011111111111111111111111111111},
{270'b111111111111111111111111111111111111100001111111111111111111111100000000011111111111111111111111000000000111111111111111111111111111111110000001111111111111000000111111111111111111100000000011111111111111000011111111111111110000011111111000011111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111}
};

localparam  int LOSE_WIDTH_X = 270;
localparam  int LOSE_HEIGHT_Y = 70;

logic [0:LOSE_HEIGHT_Y-1] [1*LOSE_WIDTH_X-1:0] lose_colors = {
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111100000111111111111111111000001111111111100000000011111111111111100001111111111111111100001111111111111111110000111111111111111111111111111110000000001111111111111111111111000000000111111111100000000000000000000000011111100001111111111111111111111111},
{270'b111111111111111111111110000011111111111111110000011111111110000000000000111111111111100001111111111111111100001111111111111111110000111111111111111111111111111000000000000011111111111111111000000000000001111111100000000000000000000000011111100001111111111111111111111111},
{270'b111111111111111111111111000011111111111111110000111111111000000000000000001111111111100001111111111111111100001111111111111111110000111111111111111111111111100000000000000000111111111111110000000000000000011111100000000000000000000000011111100001111111111111111111111111},
{270'b111111111111111111111111000001111111111111100000111111110000000000000000000111111111100001111111111111111100001111111111111111110000111111111111111111111111000000000000000000011111111111100000000000000000001111100000000000000000000000011111100001111111111111111111111111},
{270'b111111111111111111111111100000111111111111000001111111100000001111111000000011111111100001111111111111111100001111111111111111110000111111111111111111111110000000111111100000001111111111000000011111110000000111111111111110000111111111111111100001111111111111111111111111},
{270'b111111111111111111111111110000111111111111000011111111000000111111111110000001111111100001111111111111111100001111111111111111110000111111111111111111111100000011111111111000000111111111000001111111111100000111111111111110000111111111111111100001111111111111111111111111},
{270'b111111111111111111111111110000011111111110000011111110000001111111111111000000111111100001111111111111111100001111111111111111110000111111111111111111111000000111111111111100000011111110000011111111111110000011111111111110000111111111111111100001111111111111111111111111},
{270'b111111111111111111111111111000001111111100000111111110000011111111111111100000111111100001111111111111111100001111111111111111110000111111111111111111111000001111111111111110000011111110000111111111111111000011111111111110000111111111111111100001111111111111111111111111},
{270'b111111111111111111111111111100001111111100001111111100000111111111111111110000011111100001111111111111111100001111111111111111110000111111111111111111110000011111111111111111000001111110000111111111111111000011111111111110000111111111111111100001111111111111111111111111},
{270'b111111111111111111111111111100000111111000001111111100001111111111111111111000011111100001111111111111111100001111111111111111110000111111111111111111110000111111111111111111100001111110000111111111111111111111111111111110000111111111111111100001111111111111111111111111},
{270'b111111111111111111111111111110000011110000011111111100001111111111111111111000011111100001111111111111111100001111111111111111110000111111111111111111110000111111111111111111100001111110000011111111111111111111111111111110000111111111111111100001111111111111111111111111},
{270'b111111111111111111111111111111000011110000111111111000001111111111111111111000001111100001111111111111111100001111111111111111110000111111111111111111100000111111111111111111100000111111000000111111111111111111111111111110000111111111111111100001111111111111111111111111},
{270'b111111111111111111111111111111000001100000111111111000011111111111111111111100001111100001111111111111111100001111111111111111110000111111111111111111100001111111111111111111110000111111000000000111111111111111111111111110000111111111111111100001111111111111111111111111},
{270'b111111111111111111111111111111100000000001111111111000011111111111111111111100001111100001111111111111111100001111111111111111110000111111111111111111100001111111111111111111110000111111100000000000011111111111111111111110000111111111111111100001111111111111111111111111},
{270'b111111111111111111111111111111110000000011111111111000011111111111111111111100001111100001111111111111111100001111111111111111110000111111111111111111100001111111111111111111110000111111111000000000000001111111111111111110000111111111111111100001111111111111111111111111},
{270'b111111111111111111111111111111110000000011111111111000011111111111111111111100001111100001111111111111111100001111111111111111110000111111111111111111100001111111111111111111110000111111111110000000000000011111111111111110000111111111111111100001111111111111111111111111},
{270'b111111111111111111111111111111111000000111111111111000011111111111111111111100001111100001111111111111111100001111111111111111110000111111111111111111100001111111111111111111110000111111111111111000000000001111111111111110000111111111111111100001111111111111111111111111},
{270'b111111111111111111111111111111111100001111111111111000011111111111111111111100001111100001111111111111111100001111111111111111110000111111111111111111100001111111111111111111110000111111111111111111100000000111111111111110000111111111111111110011111111111111111111111111},
{270'b111111111111111111111111111111111100001111111111111000011111111111111111111100001111100001111111111111111100001111111111111111110000111111111111111111100001111111111111111111110000111111111111111111111100000011111111111110000111111111111111110011111111111111111111111111},
{270'b111111111111111111111111111111111100001111111111111000001111111111111111111000001111100001111111111111111100001111111111111111110000111111111111111111100000111111111111111111100000111111111111111111111111000001111111111110000111111111111111110011111111111111111111111111},
{270'b111111111111111111111111111111111100001111111111111100001111111111111111111000011111100001111111111111111100001111111111111111110000111111111111111111110000111111111111111111100001111100001111111111111111100001111111111110000111111111111111110011111111111111111111111111},
{270'b111111111111111111111111111111111100001111111111111100001111111111111111111000011111100001111111111111111100001111111111111111110000111111111111111111110000111111111111111111100001111100001111111111111111100001111111111110000111111111111111110011111111111111111111111111},
{270'b111111111111111111111111111111111100001111111111111100000111111111111111110000011111100000111111111111111000001111111111111111110000111111111111111111110000011111111111111111000001111100000111111111111111100001111111111110000111111111111111110011111111111111111111111111},
{270'b111111111111111111111111111111111100001111111111111110000011111111111111100000111111110000111111111111111000011111111111111111110000111111111111111111111000001111111111111110000011111110000111111111111111100001111111111110000111111111111111110011111111111111111111111111},
{270'b111111111111111111111111111111111100001111111111111110000001111111111111000000111111110000011111111111110000011111111111111111110000111111111111111111111000000111111111111100000011111110000011111111111111000001111111111110000111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111100001111111111111111000000111111111110000001111111110000001111111111100000011111111111111111110000111111111111111111111100000011111111111000000111111110000001111111111110000011111111111110000111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111100001111111111111111100000001111111000000011111111111000000011111110000000111111111111111111110000111111111111111111111110000000111111100000001111111111000000001111111000000011111111111110000111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111100001111111111111111110000000000000000000111111111111100000000000000000001111111111111111111110000000000000000000011111111000000000000000000011111111111100000000000000000000111111111111110000111111111111111100001111111111111111111111111},
{270'b111111111111111111111111111111111100001111111111111111111000000000000000001111111111111110000000000000000011111111111111111111110000000000000000000011111111100000000000000000111111111111110000000000000000001111111111111110000111111111111111100001111111111111111111111111},
{270'b111111111111111111111111111111111100001111111111111111111110000000000000111111111111111111000000000000000111111111111111111111110000000000000000000011111111111000000000000011111111111111111100000000000000111111111111111110000111111111111111100001111111111111111111111111},
{270'b111111111111111111111111111111111100001111111111111111111111100000000011111111111111111111111000000000111111111111111111111111110000000000000000000011111111111110000000001111111111111111111111000000000011111111111111111110000111111111111111100001111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111}
};


localparam  int STRIKES_WIDTH_X = 270;
localparam  int STRIKES_HEIGHT_Y = 70;

logic [0:STRIKES_HEIGHT_Y-1] [1*STRIKES_WIDTH_X-1:0] strikes_colors = {
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111100000001111111111000000000000000000011111000000000000000011111111110001111111000111111111111100001111000000000000000000111111111110000000111111111111111111111100011111111111111111000000000000000000111111000000000000000001110000000000000000000111111111111111},
{270'b111111111110000000000011111111000000000000000000011111000000000000000000111111110001111111000111111111111000011111000000000000000000111111111000000000001111111111111111111100011111111111111111000000000000000000111111000000000000000001110000000000000000000111111111111111},
{270'b111111111100000000000000111111000000000000000000011111000000000000000000011111110001111111000111111111110000111111000000000000000000111111110000000000000011111111111111111100011111111111111111000000000000000000111111000000000000000001110000000000000000000111111111111111},
{270'b111111111000001111110000011111111111110001111111111111000111111111110000011111110001111111000111111111100001111111000111111111111111111111100000111111000001111111111111111100011111111111111111000111111111111111111111000111111111111111111111111100011111111111111111111111},
{270'b111111110000111111111000011111111111110001111111111111000111111111111100001111110001111111000111111111000011111111000111111111111111111111000011111111100001111111111111111100011111111111111111000111111111111111111111000111111111111111111111111100011111111111111111111111},
{270'b111111110001111111111100001111111111110001111111111111000111111111111110001111110001111111000111111110000111111111000111111111111111111111000111111111110000111111111111111100011111111111111111000111111111111111111111000111111111111111111111111100011111111111111111111111},
{270'b111111110001111111111110001111111111110001111111111111000111111111111110001111110001111111000111111100001111111111000111111111111111111111000111111111111000111111111111111100011111111111111111000111111111111111111111000111111111111111111111111100011111111111111111111111},
{270'b111111110001111111111110001111111111110001111111111111000111111111111110001111110001111111000111111000011111111111000111111111111111111111000111111111111000111111111111111100011111111111111111000111111111111111111111000111111111111111111111111100011111111100011111111111},
{270'b111111110000111111111111111111111111110001111111111111000111111111111100001111110001111111000111110000111111111111000111111111111111111111000011111111111111111111111111111100011111111111111111000111111111111111111111000111111111111111111111111100011111111100011111111111},
{270'b111111111000011111111111111111111111110001111111111111000111111111111100001111110001111111000111100001111111111111000111111111111111111111100001111111111111111111111111111100011111111111111111000111111111111111111111000111111111111111111111111100011111111100011111111111},
{270'b111111111000000011111111111111111111110001111111111111000111111111110000011111110001111111000111000011111111111111000111111111111111111111100000001111111111111111111111111100011111111111111111000111111111111111111111000111111111111111111111111100011111111111111111111111},
{270'b111111111100000000001111111111111111110001111111111111000000000000000000111111110001111111000110000011111111111111000000000000000001111111110000000000111111111111111111111100011111111111111111000000000000000001111111000000000000000111111111111100011111111111111111111111},
{270'b111111111111000000000001111111111111110001111111111111000000000000000001111111110001111111000100000001111111111111000000000000000001111111111100000000000111111111111111111100011111111111111111000000000000000001111111000000000000000111111111111100011111111111111111111111},
{270'b111111111111110000000000011111111111110001111111111111000000000000000111111111110001111111000000010000111111111111000000000000000001111111111111000000000001111111111111111100011111111111111111000000000000000001111111000000000000000111111111111100011111111111111111111111},
{270'b111111111111111111000000001111111111110001111111111111000111111000001111111111110001111111000000111000011111111111000111111111111111111111111111111100000000111111111111111100011111111111111111000111111111111111111111000111111111111111111111111100011111111111111111111111},
{270'b111111111111111111111000001111111111110001111111111111000111111100000111111111110001111111000001111100011111111111000111111111111111111111111111111111100000111111111111111100011111111111111111000111111111111111111111000111111111111111111111111100011111111111111111111111},
{270'b111111111111111111111110000111111111110001111111111111000111111110000111111111110001111111000011111100001111111111000111111111111111111111111111111111111000011111111111111100011111111111111111000111111111111111111111000111111111111111111111111100011111111111111111111111},
{270'b111111100011111111111111000111111111110001111111111111000111111111000011111111110001111111000111111110000111111111000111111111111111111110001111111111111100011111111111111100011111111111111111000111111111111111111111000111111111111111111111111100011111111111111111111111},
{270'b111111100011111111111111000111111111110001111111111111000111111111100001111111110001111111000111111111000011111111000111111111111111111110001111111111111100011111111111111100011111111111111111000111111111111111111111000111111111111111111111111100011111111111111111111111},
{270'b111111100001111111111111000111111111110001111111111111000111111111100001111111110001111111000111111111100011111111000111111111111111111110000111111111111100011111111111111100011111111111111111000111111111111111111111000111111111111111111111111100011111111111111111111111},
{270'b111111110001111111111110000111111111110001111111111111000111111111110000111111110001111111000111111111100001111111000111111111111111111111000111111111111000011111111111111100011111111111111111000111111111111111111111000111111111111111111111111100011111111111111111111111},
{270'b111111110000011111111100001111111111110001111111111111000111111111111000011111110001111111000111111111110000111111000111111111111111111111000001111111110000111111111111111100011111111111111111000111111111111111111111000111111111111111111111111100011111111111111111111111},
{270'b111111111000000111111000001111111111110001111111111111000111111111111000011111110001111111000111111111111000111111000111111111111111111111100000011111100000111111111111111100011111111111111111000111111111111111111111000111111111111111111111111100011111111111111111111111},
{270'b111111111100000000000000011111111111110001111111111111000111111111111100001111110001111111000111111111111100011111000000000000000000011111110000000000000001111111111111111100000000000000001111000000000000000000011111000111111111111111111111111100011111111100011111111111},
{270'b111111111110000000000000111111111111110001111111111111000111111111111100001111110001111111000111111111111100001111000000000000000000011111111000000000000011111111111111111100000000000000001111000000000000000000011111000111111111111111111111111100011111111100011111111111},
{270'b111111111111100000000111111111111111110001111111111111000111111111111110000111110001111111000111111111111110000111000000000000000000011111111110000000011111111111111111111100000000000000001111000000000000000000011111000111111111111111111111111100011111111100011111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111},
{270'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111}
};


/////////////////////////////////////////////////////////

// calculate pixel location and offsets

int	inTable, inWood, inHole1, inHole2, inHole3, inHole4, inHole5,
		inHole6, hole1OffsetX, hole1OffsetY, hole2OffsetX, hole2OffsetY,
		hole3OffsetX, hole3OffsetY, hole4OffsetX, hole4OffsetY, hole5OffsetX,
		hole5OffsetY, hole6OffsetX, hole6OffsetY, inMenuText, inWinText, inLoseText, inStrikesText,
		menuTextOffsetX, menuTextOffsetY, winTextOffsetX, winTextOffsetY,
		loseTextOffsetX, loseTextOffsetY, strikesTextOffsetX, strikesTextOffsetY;

assign inTable = (pixelX > topLeftTableX && pixelX < (topLeftTableX + tableWidth) &&
						pixelY > topLeftTableY && pixelY < (topLeftTableY + tableHeight));
						
assign inGreen = (pixelX > (topLeftTableX + woodWidth) && 
						pixelX < (topLeftTableX + tableWidth - woodWidth) &&
						pixelY > (topLeftTableY + woodWidth) && 
						pixelY < (topLeftTableY + tableHeight - woodWidth));
						
assign inHole1 = ((pixelX > topLeftHole1X) && 
						(pixelX < (topLeftHole1X + HOLE_WIDTH_X)) &&
						(pixelY > topLeftHole1Y) &&
						(pixelY < (topLeftHole1Y + HOLE_HEIGHT_Y)));
						
assign hole1OffsetX = pixelX - topLeftHole1X;
assign hole1OffsetY = pixelY - topLeftHole1Y;
											
assign inHole2 = ((pixelX > topLeftHole2X) && 
						(pixelX < (topLeftHole2X + HOLE_WIDTH_X)) &&
						(pixelY > topLeftHole2Y) &&
						(pixelY < (topLeftHole2Y + HOLE_HEIGHT_Y)));
						
assign hole2OffsetX = pixelX - topLeftHole2X;
assign hole2OffsetY = pixelY - topLeftHole2Y;
						
assign inHole3 = ((pixelX > topLeftHole3X) && 
						(pixelX < (topLeftHole3X + HOLE_WIDTH_X)) &&
						(pixelY > topLeftHole3Y) &&
						(pixelY < (topLeftHole3Y + HOLE_HEIGHT_Y)));	
						
assign hole3OffsetX = pixelX - topLeftHole3X;
assign hole3OffsetY = pixelY - topLeftHole3Y;
						
assign inHole4 = ((pixelX > topLeftHole4X) && 
						(pixelX < (topLeftHole4X + HOLE_WIDTH_X)) &&
						(pixelY > topLeftHole4Y) &&
						(pixelY < (topLeftHole4Y + HOLE_HEIGHT_Y)));
						
assign hole4OffsetX = pixelX - topLeftHole4X;
assign hole4OffsetY = pixelY - topLeftHole4Y;
						
assign inHole5 = ((pixelX > topLeftHole5X) && 
						(pixelX < (topLeftHole5X + HOLE_WIDTH_X)) &&
						(pixelY > topLeftHole5Y) &&
						(pixelY < (topLeftHole5Y + HOLE_HEIGHT_Y)));	
						
assign hole5OffsetX = pixelX - topLeftHole5X;
assign hole5OffsetY = pixelY - topLeftHole5Y;
						
assign inHole6 = ((pixelX > topLeftHole6X) && 
						(pixelX < (topLeftHole6X + HOLE_WIDTH_X)) &&
						(pixelY > topLeftHole6Y) &&
						(pixelY < (topLeftHole6Y + HOLE_HEIGHT_Y)));
						
assign hole6OffsetX = pixelX - topLeftHole6X;
assign hole6OffsetY = pixelY - topLeftHole6Y;

assign inMenuText = ((pixelX > topLeftMenuX) && 
						(pixelX < (topLeftMenuX + MENU_WIDTH_X)) &&
						(pixelY > topLeftMenuY) &&
						(pixelY < (topLeftMenuY + MENU_HEIGHT_Y)));	
						
assign menuTextOffsetX = MENU_WIDTH_X - pixelX + topLeftMenuX;
assign menuTextOffsetY = pixelY - topLeftMenuY;

assign inWinText = ((pixelX > topLeftWinX) && 
						(pixelX < (topLeftWinX + WIN_WIDTH_X)) &&
						(pixelY > topLeftWinY) &&
						(pixelY < (topLeftWinY + WIN_HEIGHT_Y)));	
						
assign winTextOffsetX = WIN_WIDTH_X - pixelX + topLeftWinX;
assign winTextOffsetY = pixelY - topLeftWinY;

assign inLoseText = ((pixelX > topLeftLoseX) && 
						(pixelX < (topLeftLoseX + LOSE_WIDTH_X)) &&
						(pixelY > topLeftLoseY) &&
						(pixelY < (topLeftLoseY + LOSE_HEIGHT_Y)));	
						
assign loseTextOffsetX = LOSE_WIDTH_X - pixelX + topLeftLoseX;
assign loseTextOffsetY = pixelY - topLeftLoseY;

assign inStrikesText = ((pixelX > topLeftStrikesX) && 
						(pixelX < (topLeftStrikesX + STRIKES_WIDTH_X)) &&
						(pixelY > topLeftStrikesY) &&
						(pixelY < (topLeftStrikesY + STRIKES_HEIGHT_Y)));	
						
assign strikesTextOffsetX = STRIKES_WIDTH_X - pixelX + topLeftStrikesX;
assign strikesTextOffsetY = pixelY - topLeftStrikesY;
						
/////////////////////////////////////////////////


logic [2:0] redBits;
logic [2:0] greenBits;
logic [1:0] blueBits;

localparam logic [2:0] DARK_COLOR = 3'b111 ;// bitmap of a dark color
localparam logic [2:0] LIGHT_COLOR = 3'b000 ;// bitmap of a light color

assign BG_RGB =  {redBits , greenBits , blueBits} ; //collect color nibbles to an 8 bit word 

//----------------------------------------------------------------------------------------------
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
				redBits <= DARK_COLOR ;	
				greenBits <= DARK_COLOR  ;	
				blueBits <= DARK_COLOR ;	 
	end 
	else begin
	
	// defaults 
		greenBits <= DARK_COLOR; 
		redBits <= DARK_COLOR;
		blueBits <= DARK_COLOR;
		
		if ( inTable ) begin
			if ( inHole1 && hole_colors[hole1OffsetY][hole1OffsetX] == 1'b0 ) begin
				redBits <= LIGHT_COLOR ;	
				greenBits <= LIGHT_COLOR  ;	
				blueBits <= LIGHT_COLOR ;	
			end else if ( inHole2 && 
								hole_colors[hole2OffsetY][hole2OffsetX] == 1'b0 ) begin
				redBits <= LIGHT_COLOR ;	
				greenBits <= LIGHT_COLOR  ;	
				blueBits <= LIGHT_COLOR ;	
			end else if ( inHole3 && 
								hole_colors[hole3OffsetY][hole3OffsetX] == 1'b0 ) begin
				redBits <= LIGHT_COLOR ;	
				greenBits <= LIGHT_COLOR  ;	
				blueBits <= LIGHT_COLOR ;	
			end else if ( inHole4 && 
								hole_colors[hole4OffsetY][hole4OffsetX] == 1'b0 ) begin
				redBits <= LIGHT_COLOR ;	
				greenBits <= LIGHT_COLOR  ;	
				blueBits <= LIGHT_COLOR ;	
			end else if ( inHole5 && 
								hole_colors[hole5OffsetY][hole5OffsetX] == 1'b0 ) begin
				redBits <= LIGHT_COLOR ;	
				greenBits <= LIGHT_COLOR  ;	
				blueBits <= LIGHT_COLOR ;	
			end else if ( inHole6 && 
								hole_colors[hole6OffsetY][hole6OffsetX] == 1'b0 ) begin
				redBits <= LIGHT_COLOR ;	
				greenBits <= LIGHT_COLOR  ;	
				blueBits <= LIGHT_COLOR ;	
			end else if ( inGreen ) begin
				greenBits <= 3'b100; 
				redBits <= 3'b000;
				blueBits <= 2'b00;
			end else begin //in edge
				greenBits <= 3'b100; 
				redBits <= 3'b100;
				blueBits <= 2'b01;
			end
		end
		
		if (menu_state == 1'b1 && inMenuText &&
			 menu_colors[menuTextOffsetY][menuTextOffsetX] == 1'b0) begin
				redBits <= LIGHT_COLOR ;	
				greenBits <= LIGHT_COLOR  ;	
				blueBits <= LIGHT_COLOR ;	 
		end
		
		if (end_state == 1'b1 && win == 1'b1 && inWinText &&
			 win_colors[winTextOffsetY][winTextOffsetX] == 1'b0) begin
				redBits <= LIGHT_COLOR ;	
				greenBits <= LIGHT_COLOR  ;	
				blueBits <= LIGHT_COLOR ; 
		end
		
		if (end_state == 1'b1 && win == 1'b0 && inLoseText &&
			 lose_colors[loseTextOffsetY][loseTextOffsetX] == 1'b0) begin
				redBits <= LIGHT_COLOR ;	
				greenBits <= LIGHT_COLOR  ;	
				blueBits <= LIGHT_COLOR ;
		end	

		if (inStrikesText && strikes_colors[strikesTextOffsetY][strikesTextOffsetX] == 1'b0) begin
				redBits <= LIGHT_COLOR ;	
				greenBits <= LIGHT_COLOR  ;	
				blueBits <= LIGHT_COLOR ;
		end		


		
	end; 	
end 

endmodule
