// (c) Technion IIT, Department of Electrical Engineering 2019 
// Written By Natan Kaminsky and Nimrod Barazani June 2019

module stick_move 	
 ( 
   input	   logic  clk,
	input	   logic  resetN, 
	input	   logic  startOfFrame,
	input	   logic  up_pressed,
	input	   logic  down_pressed,
	input	   logic  space_pressed,
	input	   logic  game_state,
	input	   logic  no_moving_flag,
	input	   logic  [10:0] whiteBallTopLeftX,
	input	   logic  [10:0] whiteBallTopLeftY,
	output   logic  [10:0] stickCenterX,
	output   logic  [10:0] stickCenterY,
   output   int velocityX,
	output   int velocityY,
	output   logic  [9:0] angle
	 
  ) ;

localparam int MAX_ANGLE = 359;
const logic [0:MAX_ANGLE] [15:0] sin_table = {16'h0000,16'h0008,16'h0011,16'h001A,16'h0023,16'h002C,16'h0035,16'h003E,16'h0047,16'h0050,16'h0058,16'h0061,
16'h006A,16'h0073,16'h007B,16'h0084,16'h008D,16'h0095,16'h009E,16'h00A6,16'h00AF,16'h00B7,16'h00BF,16'h00C8,16'h00D0,16'h00D8,16'h00E0,16'h00E8,16'h00F0,
16'h00F8,16'h00FF,16'h0107,16'h010F,16'h0116,16'h011E,16'h0125,16'h012C,16'h0134,16'h013B,16'h0142,16'h0149,16'h014F,16'h0156,16'h015D,16'h0163,16'h016A,
16'h0170,16'h0176,16'h017C,16'h0182,16'h0188,16'h018D,16'h0193,16'h0198,16'h019E,16'h01A3,16'h01A8,16'h01AD,16'h01B2,16'h01B6,16'h01BB,16'h01BF,16'h01C4,
16'h01C8,16'h01CC,16'h01D0,16'h01D3,16'h01D7,16'h01DA,16'h01DD,16'h01E1,16'h01E4,16'h01E6,16'h01E9,16'h01EC,16'h01EE,16'h01F0,16'h01F2,16'h01F4,16'h01F6,
16'h01F8,16'h01F9,16'h01FB,16'h01FC,16'h01FD,16'h01FE,16'h01FE,16'h01FF,16'h01FF,16'h01FF,16'h0200,16'h01FF,16'h01FF,16'h01FF,16'h01FE,16'h01FE,16'h01FD,
16'h01FC,16'h01FB,16'h01F9,16'h01F8,16'h01F6,16'h01F4,16'h01F2,16'h01F0,16'h01EE,16'h01EC,16'h01E9,16'h01E6,16'h01E4,16'h01E1,16'h01DD,16'h01DA,16'h01D7,
16'h01D3,16'h01D0,16'h01CC,16'h01C8,16'h01C4,16'h01BF,16'h01BB,16'h01B6,16'h01B2,16'h01AD,16'h01A8,16'h01A3,16'h019E,16'h0198,16'h0193,16'h018D,16'h0188,
16'h0182,16'h017C,16'h0176,16'h0170,16'h016A,16'h0163,16'h015D,16'h0156,16'h014F,16'h0149,16'h0142,16'h013B,16'h0134,16'h012C,16'h0125,16'h011E,16'h0116,
16'h010F,16'h0107,16'h00FF,16'h00F8,16'h00F0,16'h00E8,16'h00E0,16'h00D8,16'h00D0,16'h00C8,16'h00BF,16'h00B7,16'h00AF,16'h00A6,16'h009E,16'h0095,16'h008D,
16'h0084,16'h007B,16'h0073,16'h006A,16'h0061,16'h0058,16'h0050,16'h0047,16'h003E,16'h0035,16'h002C,16'h0023,16'h001A,16'h0011,16'h0008,16'h0000,16'hFFF8,
16'hFFEF,16'hFFE6,16'hFFDD,16'hFFD4,16'hFFCB,16'hFFC2,16'hFFB9,16'hFFB0,16'hFFA8,16'hFF9F,16'hFF96,16'hFF8D,16'hFF85,16'hFF7C,16'hFF73,16'hFF6B,16'hFF62,
16'hFF5A,16'hFF51,16'hFF49,16'hFF41,16'hFF38,16'hFF30,16'hFF28,16'hFF20,16'hFF18,16'hFF10,16'hFF08,16'hFF00,16'hFEF9,16'hFEF1,16'hFEEA,16'hFEE2,16'hFEDB,
16'hFED4,16'hFECC,16'hFEC5,16'hFEBE,16'hFEB7,16'hFEB1,16'hFEAA,16'hFEA3,16'hFE9D,16'hFE96,16'hFE90,16'hFE8A,16'hFE84,16'hFE7E,16'hFE78,16'hFE73,16'hFE6D,
16'hFE68,16'hFE62,16'hFE5D,16'hFE58,16'hFE53,16'hFE4E,16'hFE4A,16'hFE45,16'hFE41,16'hFE3C,16'hFE38,16'hFE34,16'hFE30,16'hFE2D,16'hFE29,16'hFE26,16'hFE23,
16'hFE1F,16'hFE1C,16'hFE1A,16'hFE17,16'hFE14,16'hFE12,16'hFE10,16'hFE0E,16'hFE0C,16'hFE0A,16'hFE08,16'hFE07,16'hFE05,16'hFE04,16'hFE03,16'hFE02,16'hFE02,
16'hFE01,16'hFE01,16'hFE01,16'hFE00,16'hFE01,16'hFE01,16'hFE01,16'hFE02,16'hFE02,16'hFE03,16'hFE04,16'hFE05,16'hFE07,16'hFE08,16'hFE0A,16'hFE0C,16'hFE0E,
16'hFE10,16'hFE12,16'hFE14,16'hFE17,16'hFE1A,16'hFE1C,16'hFE1F,16'hFE23,16'hFE26,16'hFE29,16'hFE2D,16'hFE30,16'hFE34,16'hFE38,16'hFE3C,16'hFE41,16'hFE45,
16'hFE4A,16'hFE4E,16'hFE53,16'hFE58,16'hFE5D,16'hFE62,16'hFE68,16'hFE6D,16'hFE73,16'hFE78,16'hFE7E,16'hFE84,16'hFE8A,16'hFE90,16'hFE96,16'hFE9D,16'hFEA3,
16'hFEAA,16'hFEB1,16'hFEB7,16'hFEBE,16'hFEC5,16'hFECC,16'hFED4,16'hFEDB,16'hFEE2,16'hFEEA,16'hFEF1,16'hFEF9,16'hFF00,16'hFF08,16'hFF10,16'hFF18,16'hFF20,
16'hFF28,16'hFF30,16'hFF38,16'hFF41,16'hFF49,16'hFF51,16'hFF5A,16'hFF62,16'hFF6B,16'hFF73,16'hFF7C,16'hFF85,16'hFF8D,16'hFF96,16'hFF9F,16'hFFA8,16'hFFB0,
16'hFFB9,16'hFFC2,16'hFFCB,16'hFFD4,16'hFFDD,16'hFFE6,16'hFFEF,16'hFFF8  };
 
 const logic [0:MAX_ANGLE] [15:0] cos_table = {16'h0200,16'h01FF,16'h01FF,16'h01FF,16'h01FE,16'h01FE,16'h01FD,16'h01FC,16'h01FB,16'h01F9,16'h01F8,16'h01F6,
16'h01F4,16'h01F2,16'h01F0,16'h01EE,16'h01EC,16'h01E9,16'h01E6,16'h01E4,16'h01E1,16'h01DD,16'h01DA,16'h01D7,16'h01D3,16'h01D0,16'h01CC,16'h01C8,16'h01C4,
16'h01BF,16'h01BB,16'h01B6,16'h01B2,16'h01AD,16'h01A8,16'h01A3,16'h019E,16'h0198,16'h0193,16'h018D,16'h0188,16'h0182,16'h017C,16'h0176,16'h0170,16'h016A,
16'h0163,16'h015D,16'h0156,16'h014F,16'h0149,16'h0142,16'h013B,16'h0134,16'h012C,16'h0125,16'h011E,16'h0116,16'h010F,16'h0107,16'h0100,16'h00F8,16'h00F0,
16'h00E8,16'h00E0,16'h00D8,16'h00D0,16'h00C8,16'h00BF,16'h00B7,16'h00AF,16'h00A6,16'h009E,16'h0095,16'h008D,16'h0084,16'h007B,16'h0073,16'h006A,16'h0061,
16'h0058,16'h0050,16'h0047,16'h003E,16'h0035,16'h002C,16'h0023,16'h001A,16'h0011,16'h0008,16'h0000,16'hFFF8,16'hFFEF,16'hFFE6,16'hFFDD,16'hFFD4,16'hFFCB,
16'hFFC2,16'hFFB9,16'hFFB0,16'hFFA8,16'hFF9F,16'hFF96,16'hFF8D,16'hFF85,16'hFF7C,16'hFF73,16'hFF6B,16'hFF62,16'hFF5A,16'hFF51,16'hFF49,16'hFF41,16'hFF38,
16'hFF30,16'hFF28,16'hFF20,16'hFF18,16'hFF10,16'hFF08,16'hFF01,16'hFEF9,16'hFEF1,16'hFEEA,16'hFEE2,16'hFEDB,16'hFED4,16'hFECC,16'hFEC5,16'hFEBE,16'hFEB7,
16'hFEB1,16'hFEAA,16'hFEA3,16'hFE9D,16'hFE96,16'hFE90,16'hFE8A,16'hFE84,16'hFE7E,16'hFE78,16'hFE73,16'hFE6D,16'hFE68,16'hFE62,16'hFE5D,16'hFE58,16'hFE53,
16'hFE4E,16'hFE4A,16'hFE45,16'hFE41,16'hFE3C,16'hFE38,16'hFE34,16'hFE30,16'hFE2D,16'hFE29,16'hFE26,16'hFE23,16'hFE1F,16'hFE1C,16'hFE1A,16'hFE17,16'hFE14,
16'hFE12,16'hFE10,16'hFE0E,16'hFE0C,16'hFE0A,16'hFE08,16'hFE07,16'hFE05,16'hFE04,16'hFE03,16'hFE02,16'hFE02,16'hFE01,16'hFE01,16'hFE01,16'hFE00,16'hFE01,
16'hFE01,16'hFE01,16'hFE02,16'hFE02,16'hFE03,16'hFE04,16'hFE05,16'hFE07,16'hFE08,16'hFE0A,16'hFE0C,16'hFE0E,16'hFE10,16'hFE12,16'hFE14,16'hFE17,16'hFE1A,
16'hFE1C,16'hFE1F,16'hFE23,16'hFE26,16'hFE29,16'hFE2D,16'hFE30,16'hFE34,16'hFE38,16'hFE3C,16'hFE41,16'hFE45,16'hFE4A,16'hFE4E,16'hFE53,16'hFE58,16'hFE5D,
16'hFE62,16'hFE68,16'hFE6D,16'hFE73,16'hFE78,16'hFE7E,16'hFE84,16'hFE8A,16'hFE90,16'hFE96,16'hFE9D,16'hFEA3,16'hFEAA,16'hFEB1,16'hFEB7,16'hFEBE,16'hFEC5,
16'hFECC,16'hFED4,16'hFEDB,16'hFEE2,16'hFEEA,16'hFEF1,16'hFEF9,16'hFF00,16'hFF08,16'hFF10,16'hFF18,16'hFF20,16'hFF28,16'hFF30,16'hFF38,16'hFF41,16'hFF49,
16'hFF51,16'hFF5A,16'hFF62,16'hFF6B,16'hFF73,16'hFF7C,16'hFF85,16'hFF8D,16'hFF96,16'hFF9F,16'hFFA8,16'hFFB0,16'hFFB9,16'hFFC2,16'hFFCB,16'hFFD4,16'hFFDD,
16'hFFE6,16'hFFEF,16'hFFF8,16'h0000,16'h0008,16'h0011,16'h001A,16'h0023,16'h002C,16'h0035,16'h003E,16'h0047,16'h0050,16'h0058,16'h0061,16'h006A,16'h0073,
16'h007B,16'h0084,16'h008D,16'h0095,16'h009E,16'h00A6,16'h00AF,16'h00B7,16'h00BF,16'h00C8,16'h00D0,16'h00D8,16'h00E0,16'h00E8,16'h00F0,16'h00F8,16'h0100,
16'h0107,16'h010F,16'h0116,16'h011E,16'h0125,16'h012C,16'h0134,16'h013B,16'h0142,16'h0149,16'h014F,16'h0156,16'h015D,16'h0163,16'h016A,16'h0170,16'h0176,
16'h017C,16'h0182,16'h0188,16'h018D,16'h0193,16'h0198,16'h019E,16'h01A3,16'h01A8,16'h01AD,16'h01B2,16'h01B6,16'h01BB,16'h01BF,16'h01C4,16'h01C8,16'h01CC,
16'h01D0,16'h01D3,16'h01D7,16'h01DA,16'h01DD,16'h01E1,16'h01E4,16'h01E6,16'h01E9,16'h01EC,16'h01EE,16'h01F0,16'h01F2,16'h01F4,16'h01F6,16'h01F8,16'h01F9,
16'h01FB,16'h01FC,16'h01FD,16'h01FE,16'h01FE,16'h01FF,16'h01FF,16'h01FF };
    

parameter int INITIAL_X = 320; //TBD
parameter int INITIAL_Y = 240; //TBD
parameter int INITIAL_VELOCITY = 10; //TBD
parameter int MAX_VELOCITY = 510;
 
int BALLWIDTH = 16;
int BALLHEIGHT = 16;

int VELOCITY_ABS = 5; //TBD
int velX_temp;
int velY_temp;
int SIN,COS;

assign SIN = {{16{sin_table[angle][15]}},sin_table[angle]};
assign COS = {{16{cos_table[angle][15]}},cos_table[angle]};

	 
	 


//position calculate
always_ff @(posedge clk or negedge resetN) begin
if(!resetN)
	begin
		stickCenterX	<= INITIAL_X + BALLWIDTH/2;
		stickCenterY	<= INITIAL_Y + BALLHEIGHT/2;
	end
	else begin
			stickCenterX  	<= whiteBallTopLeftX + BALLWIDTH/2;
			stickCenterY	<= whiteBallTopLeftY + BALLHEIGHT/2;
	end
	 
end // end always_ff position calculate


//angle calculation
always_ff @(posedge clk or negedge resetN) begin
	if(!resetN)
		angle	<= 0;
		
	else if (startOfFrame == 1'b1) begin
		if (no_moving_flag == 1'b0 || game_state == 1'b0) 
			angle	<= 0;
		else begin
			if (up_pressed == 1'b1) begin
				if (angle == MAX_ANGLE)
					angle <= 0;
				else
					angle++;
			end//end if up_pressed
			
			else if (down_pressed == 1'b1) begin
				if (angle == 0)
					angle <= MAX_ANGLE;
				else
					angle--;
			end//end if down_pressed
		end
		
	end
	 
end // end always_ff angle calculate


//VELOCITY calculation
always_ff @(posedge clk or negedge resetN) begin
	if(!resetN)
		VELOCITY_ABS	<= INITIAL_VELOCITY;
	else if (startOfFrame == 1'b1) begin
		
		if (no_moving_flag == 1'b0 || game_state == 1'b0) begin
			VELOCITY_ABS	<= INITIAL_VELOCITY;
		end//end if there is a moving ball
		
		else if (space_pressed == 1'b1) begin
			if (VELOCITY_ABS < MAX_VELOCITY)
				VELOCITY_ABS<=VELOCITY_ABS+5;
		end
		
	end
	 
end // end always_ff VELOCITY calculate
 
 

   
	
	
	
	
	
 
// combinational part 

assign	velocityX = (VELOCITY_ABS*COS)/512;
assign	velocityY = (VELOCITY_ABS*SIN)/512; 
	
 
endmodule

